library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_TMR is
end tb_TMR;

architecture Behavioral of tb_TMR is
    constant CLK_PERIOD : time := 1.55 ns;
    
    signal clk : std_logic := '0';
    signal rst : std_logic := '0';
    signal ce : std_logic := '0';
    signal A : std_logic_vector(7 downto 0) := (others => '0');
    signal B : std_logic_vector(7 downto 0) := (others => '0');
    signal OP : std_logic_vector(2 downto 0) := (others => '0');
    signal flag : std_logic;
    signal result : std_logic_vector(7 downto 0);
begin
    uut : entity work.TMR
        port map(
            clk => clk,
            rst => rst,
            ce => ce,
            A => A,
            B => B,
            OP => OP,
            flag => flag,
            result => result         
        );
    
    clk_process : process
    begin
        while true loop
           clk <= '0';
           wait for CLK_PERIOD;
           clk <= '1';
           wait for CLK_PERIOD;
        end loop;
    end process;    
    
    stim_process : process
    begin
        ce <= '0';
        rst <= '1';
        wait until rising_edge(clk);
        rst <= '0';
        ce <= '1'; 
        
        A <= std_logic_vector(to_signed(1,8));
        B <= std_logic_vector(to_signed(2,8));
        OP <= "000";
        
        wait until rising_edge(clk);
 
        A <= std_logic_vector(to_signed(2,8));
        B <= std_logic_vector(to_signed(1,8));
        OP <= "001";
        
        wait until rising_edge(clk);
        
        A <= std_logic_vector(to_signed(5,8));
        B <= std_logic_vector(to_signed(3,8));
        OP <= "001";
        
        wait until rising_edge(clk);
        
        wait;
    end process;
end Behavioral;
